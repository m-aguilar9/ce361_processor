`timescale 1ns/10ps

module not_gate (x, z);
  input x;
  output z;
  
  assign z = ~x ;
  
  
endmodule
  




